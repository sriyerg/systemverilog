module top;

  foo u_foo();

endmodule
