config ip_cfg;
  design dv.foo_tb;
  default liblist ip dv work;
endconfig
