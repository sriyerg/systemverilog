config foundry_cfg;
  design dv.top_tb;
  default liblist foundry system ip dv work;
endconfig
