config system_cfg;
  design dv.top_tb;
  default liblist system ip dv work;
endconfig
